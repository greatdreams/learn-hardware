// ????????
module my_nor(out, a,b);
output out;
input a, b;

//internal wires
wire c;

//??????
supply1 pwr;   // pwr???Vdd
supply0 gnd;  // gnd???Vss(?)


// ????PMOS??
pmos (c, pwr, b);
pmos (out, c, a);

// ????NMOS??
nmos(out, gnd, a);
nmos(out, gnd, b);



endmodule