// ?????????????
module my_mux(out, s, i0, i1);

output out;
input s, i0, i1;

// ????
wire sbar; // s??
// ??s??

// ????????CMOS??
my_nor nt(sbar, s, s);

// ??(????)CMOS??
cmos(out, i0, sbar, s);
cmos (out, i1, s, sbar);

endmodule